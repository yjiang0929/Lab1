`define AND and #30
`define OR or #30
`define NOT not #10

module structuralAnd
(
    output[31:0] out,
    input[31:0] A,
    input[31:0] B
);


`AND and0(out[0],A[0],B[0]);
`AND and1(out[1],A[1],B[1]);
`AND and2(out[2],A[2],B[2]);
`AND and3(out[3],A[3],B[3]);
`AND and4(out[4],A[4],B[4]);
`AND and5(out[5],A[5],B[5]);
`AND and6(out[6],A[6],B[6]);
`AND and7(out[7],A[7],B[7]);
`AND and8(out[8],A[8],B[8]);
`AND and9(out[9],A[9],B[9]);
`AND and10(out[10],A[10],B[10]);
`AND and11(out[11],A[11],B[11]);
`AND and12(out[12],A[12],B[12]);
`AND and13(out[13],A[13],B[13]);
`AND and14(out[14],A[14],B[14]);
`AND and15(out[15],A[15],B[15]);
`AND and16(out[16],A[16],B[16]);
`AND and17(out[17],A[17],B[17]);
`AND and18(out[18],A[18],B[18]);
`AND and19(out[19],A[19],B[19]);
`AND and20(out[20],A[20],B[20]);
`AND and21(out[21],A[21],B[21]);
`AND and22(out[22],A[22],B[22]);
`AND and23(out[23],A[23],B[23]);
`AND and24(out[24],A[24],B[24]);
`AND and25(out[25],A[25],B[25]);
`AND and26(out[26],A[26],B[26]);
`AND and27(out[27],A[27],B[27]);
`AND and28(out[28],A[28],B[28]);
`AND and29(out[29],A[29],B[29]);
`AND and30(out[30],A[30],B[30]);
`AND and31(out[31],A[31],B[31]);


endmodule
